`timescale 1ns / 1ps

module intc(
    input iack,
    input [3:0] done,
    output irq,
    output addr
    );
    
    // TODO Add priority selection
    
endmodule
